entity Mandelbrot_tb is
end Mandelbrot_tb;

architecture sim of Mandelbrot_tb is
begin
end sim;